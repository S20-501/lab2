	-- megafunction wizard: %FIFO%
	-- GENERATION: STANDARD
	-- VERSION: WM1.0
	-- MODULE: scfifo 

	-- ============================================================
	-- File Name: fifoWithrst.vhd
	-- Megafunction Name(s):
	-- 			scfifo
	--
	-- Simulation Library Files(s):
	-- 			altera_mf
	-- ============================================================
	-- ************************************************************
	-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
	--
	-- 18.0.0 Build 614 04/24/2018 SJ Standard Edition
	-- ************************************************************


	--Copyright (C) 2018  Intel Corporation. All rights reserved.
	--Your use of Intel Corporation's design tools, logic functions 
	--and other software and tools, and its AMPP partner logic 
	--functions, and any output files from any of the foregoing 
	--(including device programming or simulation files), and any 
	--associated documentation or information are expressly subject 
	--to the terms and conditions of the Intel Program License 
	--Subscription Agreement, the Intel Quartus Prime License Agreement,
	--the Intel FPGA IP License Agreement, or other applicable license
	--agreement, including, without limitation, that your use is for
	--the sole purpose of programming logic devices manufactured by
	--Intel and sold by Intel or its authorized distributors.  Please
	--refer to the applicable agreement for further details.


	LIBRARY ieee;
	USE ieee.std_logic_1164.all;

	LIBRARY altera_mf;
	USE altera_mf.all;

	ENTITY GSMRegistr_FIFO IS
		PORT
		(
			aclr		: IN STD_LOGIC ;
			clock		: IN STD_LOGIC ;
			data		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			rdreq		: IN STD_LOGIC ;
			wrreq		: IN STD_LOGIC ;
			almost_full		: OUT STD_LOGIC ;
			empty		: OUT STD_LOGIC ;
			q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			usedw		: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
		);
	END GSMRegistr_FIFO;


	ARCHITECTURE SYN OF gsmregistr_fifo IS

		SIGNAL sub_wire0	: STD_LOGIC ;
		SIGNAL sub_wire1	: STD_LOGIC ;
		SIGNAL sub_wire2	: STD_LOGIC_VECTOR (15 DOWNTO 0);
		SIGNAL sub_wire3	: STD_LOGIC_VECTOR (9 DOWNTO 0);



		COMPONENT scfifo
		GENERIC (
			add_ram_output_register		: STRING;
			almost_full_value		: NATURAL;
			intended_device_family		: STRING;
			lpm_numwords		: NATURAL;
			lpm_showahead		: STRING;
			lpm_type		: STRING;
			lpm_width		: NATURAL;
			lpm_widthu		: NATURAL;
			overflow_checking		: STRING;
			underflow_checking		: STRING;
			use_eab		: STRING
		);
		PORT (
				aclr	: IN STD_LOGIC ;
				clock	: IN STD_LOGIC ;
				data	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				rdreq	: IN STD_LOGIC ;
				wrreq	: IN STD_LOGIC ;
				almost_full	: OUT STD_LOGIC ;
				empty	: OUT STD_LOGIC ;
				q	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
				usedw	: OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
		);
		END COMPONENT;

	BEGIN
		almost_full    <= sub_wire0;
		empty    <= sub_wire1;
		q    <= sub_wire2(15 DOWNTO 0);
		usedw    <= sub_wire3(9 DOWNTO 0);

		scfifo_component : scfifo
		GENERIC MAP (
			add_ram_output_register => "OFF",
			almost_full_value => 1023,
			intended_device_family => "Cyclone 10 LP",
			lpm_numwords => 1024,
			lpm_showahead => "OFF",
			lpm_type => "scfifo",
			lpm_width => 16,
			lpm_widthu => 10,
			overflow_checking => "ON",
			underflow_checking => "ON",
			use_eab => "ON"
		)
		PORT MAP (
			aclr => aclr,
			clock => clock,
			data => data,
			rdreq => rdreq,
			wrreq => wrreq,
			almost_full => sub_wire0,
			empty => sub_wire1,
			q => sub_wire2,
			usedw => sub_wire3
		);



	END SYN;

	-- ============================================================
	-- CNX file retrieval info
	-- ============================================================
	-- Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
	-- Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
	-- Retrieval info: PRIVATE: AlmostFull NUMERIC "1"
	-- Retrieval info: PRIVATE: AlmostFullThr NUMERIC "1023"
	-- Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
	-- Retrieval info: PRIVATE: Clock NUMERIC "0"
	-- Retrieval info: PRIVATE: Depth NUMERIC "1024"
	-- Retrieval info: PRIVATE: Empty NUMERIC "1"
	-- Retrieval info: PRIVATE: Full NUMERIC "0"
	-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone 10 LP"
	-- Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
	-- Retrieval info: PRIVATE: LegacyRREQ NUMERIC "1"
	-- Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
	-- Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
	-- Retrieval info: PRIVATE: Optimize NUMERIC "0"
	-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
	-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
	-- Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
	-- Retrieval info: PRIVATE: UsedW NUMERIC "1"
	-- Retrieval info: PRIVATE: Width NUMERIC "16"
	-- Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
	-- Retrieval info: PRIVATE: diff_widths NUMERIC "0"
	-- Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
	-- Retrieval info: PRIVATE: output_width NUMERIC "16"
	-- Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
	-- Retrieval info: PRIVATE: rsFull NUMERIC "0"
	-- Retrieval info: PRIVATE: rsUsedW NUMERIC "0"
	-- Retrieval info: PRIVATE: sc_aclr NUMERIC "1"
	-- Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
	-- Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
	-- Retrieval info: PRIVATE: wsFull NUMERIC "1"
	-- Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
	-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
	-- Retrieval info: CONSTANT: ADD_RAM_OUTPUT_REGISTER STRING "OFF"
	-- Retrieval info: CONSTANT: ALMOST_FULL_VALUE NUMERIC "1023"
	-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone 10 LP"
	-- Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "1024"
	-- Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "OFF"
	-- Retrieval info: CONSTANT: LPM_TYPE STRING "scfifo"
	-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "16"
	-- Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "10"
	-- Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
	-- Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
	-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
	-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
	-- Retrieval info: USED_PORT: almost_full 0 0 0 0 OUTPUT NODEFVAL "almost_full"
	-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
	-- Retrieval info: USED_PORT: data 0 0 16 0 INPUT NODEFVAL "data[15..0]"
	-- Retrieval info: USED_PORT: empty 0 0 0 0 OUTPUT NODEFVAL "empty"
	-- Retrieval info: USED_PORT: q 0 0 16 0 OUTPUT NODEFVAL "q[15..0]"
	-- Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL "rdreq"
	-- Retrieval info: USED_PORT: usedw 0 0 10 0 OUTPUT NODEFVAL "usedw[9..0]"
	-- Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL "wrreq"
	-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
	-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
	-- Retrieval info: CONNECT: @data 0 0 16 0 data 0 0 16 0
	-- Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
	-- Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
	-- Retrieval info: CONNECT: almost_full 0 0 0 0 @almost_full 0 0 0 0
	-- Retrieval info: CONNECT: empty 0 0 0 0 @empty 0 0 0 0
	-- Retrieval info: CONNECT: q 0 0 16 0 @q 0 0 16 0
	-- Retrieval info: CONNECT: usedw 0 0 10 0 @usedw 0 0 10 0
	-- Retrieval info: GEN_FILE: TYPE_NORMAL fifoWithrst.vhd TRUE
	-- Retrieval info: GEN_FILE: TYPE_NORMAL fifoWithrst.inc FALSE
	-- Retrieval info: GEN_FILE: TYPE_NORMAL fifoWithrst.cmp TRUE
	-- Retrieval info: GEN_FILE: TYPE_NORMAL fifoWithrst.bsf FALSE
	-- Retrieval info: GEN_FILE: TYPE_NORMAL fifoWithrst_inst.vhd FALSE
	-- Retrieval info: LIB_FILE: altera_mf
