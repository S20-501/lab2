	library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
LIBRARY altera_mf;
USE altera_mf.all;

entity Tester is
  port (
    -- входные данные с FT
    FT2232H_FSDI : in std_logic;
    -- Входной тактовый сигнал для микросхемы FT2232H
    FT2232H_FSCLK : in std_logic;
    -- общие сигналы
    tester_clk : out std_logic := '0';
    tester_reset : out std_logic := '1';
    -- готовность FT к приму данных (0)
    FT2232H_FSCTS : out std_logic := '1';
    -- канал передачи данных к FT
    FT2232H_FSDO : out std_logic := '1'
  );
end Tester;


-- симуляция побитовой оптравки данных
architecture tester_top of Tester is
  --общее...
  constant TbPeriod : time := 2 ps;
  signal TbClock : std_logic := '1';
  signal TbSimEnded : std_logic := '0';
  --увеличивающийся при каждом запросе TID
  signal TID_count : std_logic_vector(7 downto 0) := "00000000";
  --увеличивающийся при записи FT2232H_FSDI счетчик
  signal FSDI_count : std_logic_vector(3 downto 0) := "0000";
  --активен(1), если в данный момент идет запись в CTS
  signal CTS_open_r : std_logic := '0';
  --нужен для просмотра отправляемой информации
  signal test_FullHeader : std_logic_vector(47 downto 0);
  --проверка конкатенации с выводом результата


  function Test_Concatination(
    constant BCount : in std_logic_vector(9 downto 0);
    constant FB : in std_logic;
    constant Cmd : in std_logic_vector(2 downto 0);
    constant TID_count : in std_logic_vector(7 downto 0);
    constant Addr : in std_logic_vector(15 downto 0)
  ) return std_logic_vector is
    variable FullHeader : std_logic_vector(47 downto 0);
  begin

    FullHeader := BCount & "00" & FB & Cmd & "00000000" & TID_count & Addr;
    --FullHeader := Addr & "00000000" & TID_count & BCount & "00" & FB & Cmd;
    return FullHeader;

  end function Test_Concatination;


  procedure skiptime(time_count : in integer) is
  begin

    count_time : for k in 0 to time_count - 1 loop
      wait until rising_edge(TbClock);
    end loop count_time;

  end;


  --увеличение счетчика запросов
  function RecalculationTID(TID_count : in std_logic_vector(7 downto 0)) return std_logic_vector is
    variable result : std_logic_vector(7 downto 0);
  begin

    if TID_count = "11111111" then
      result := "00000000";
    else
      result := std_logic_vector(to_unsigned(to_integer(unsigned(TID_count)) + 1, 8));
    end if;
    return result;

  end function RecalculationTID;


  --процедура записи
  procedure WriteCommand(
    -- количество байт данных
    constant BCount : in std_logic_vector(9 downto 0);
    -- FeedBack наличие 1 - необходимость отправки на  хост для подтверждения приема и корректного анализа
    constant FB : in std_logic;
    -- команда
    constant Cmd : in std_logic_vector(2 downto 0);
    -- идентификатор транзакции
    constant TID_count : in std_logic_vector(7 downto 0);
    -- Адрес назначения (источника) данных
    constant Addr : in std_logic_vector(15 downto 0);
    --данные для записи
    constant data : in std_logic_vector;
    --выходы для записи
    signal FT2232H_FSDO : out std_logic
  )is
    variable FullHeader : std_logic_vector(0 to 47);
  begin

    FullHeader := Addr & "00000000" & TID_count & BCount & "00" & FB & Cmd;

    --циклическая запись заголовка
    full_write : for k in 0 to 5 loop
      -- запись Start bit (==0), если 1 то ошибка
      if (k /= 0) then
        wait until rising_edge(TbClock);
      end if;
      FT2232H_FSDO <= '0';
      --запись 8 значащих бит
      write8bit : for i in 0 to 7 loop
        wait until rising_edge(TbClock);
        --FT2232H_FSDO <= FullHeader(i + k*8);
        FT2232H_FSDO <= FullHeader(47 - (k * 8 + i));--записываемый бит
      end loop write8bit;
      -- запись Source bit
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '1';
    end loop full_write;

    if (BCount(0) /= '1') then
      --циклическая запись данных
      data_write1 : for g in 0 to ((to_integer(unsigned(BCount)))/2 - 1) loop
        -- запись Start bit (==0), если 1 то ошибка
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= '0';
        --запись 16 значащих бит
        write16bit_data1 : for n in 15 downto 0 loop
          if (n = 7) then
            wait until rising_edge(TbClock);
            FT2232H_FSDO <= '1';
            wait until rising_edge(TbClock);
            FT2232H_FSDO <= '0';
          end if;

          wait until rising_edge(TbClock);
          FT2232H_FSDO <= data(n + g * 16);
        end loop write16bit_data1;
        -- запись Source bit
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= '1';
      end loop data_write1;

    else

	 
	 --циклическая запись данных
      data_write2 : for g in 0 to ((to_integer(unsigned(BCount)))/2 - 1) loop
        -- запись Start bit (==0), если 1 то ошибка
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= '0';
        --запись 16 значащих бит
        write16bit_data2 : for n in 15 downto 0 loop
          if (n = 7) then
            wait until rising_edge(TbClock);
            FT2232H_FSDO <= '1';
            wait until rising_edge(TbClock);
            FT2232H_FSDO <= '0';
          end if;

          wait until rising_edge(TbClock);
          FT2232H_FSDO <= data(n + g * 16);
        end loop write16bit_data2;
        -- запись Source bit
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= '1';
      end loop data_write2;
	 
	 
      --значащая наоборот, а потом нули
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '0';
      write8bit_data1 : for q in ((to_integer(unsigned(BCount)))*8-1) downto ((to_integer(unsigned(BCount)))*8-8) loop
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= data(q);
      end loop write8bit_data1;
		
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '1';
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '0';
		
      write8bit_data2 : for q in 7 downto 0 loop
        wait until rising_edge(TbClock);
        FT2232H_FSDO <= '0';
      end loop write8bit_data2;
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '1';

    end if;

  end procedure WriteCommand;
  --процедура чтения
  procedure ReadCommand(
    -- количество байт данных
    constant BCount : in std_logic_vector(9 downto 0);
    -- FeedBack наличие 1 - необходимость отправки на  хост для подтверждения приема и корректного анализа
    constant FB : in std_logic;
    -- команда
    constant Cmd : in std_logic_vector(2 downto 0);
    -- идентификатор транзакции
    constant TID_couunt : in std_logic_vector(7 downto 0);
    -- Адрес назначения (источника) данных
    constant Addr : in std_logic_vector(15 downto 0);
    signal FT2232H_FSDO : out std_logic
  )is
    variable FullHeader : std_logic_vector(0 to 47);
  begin

    FullHeader := Addr & "00000000" & TID_count & BCount & "00" & FB & Cmd; 

    --циклическая запись заголовка
    full_write : for k in 0 to 5 loop
      -- запись Start bit (==0), если 1 то ошибка
      if (k /= 0) then
        wait until rising_edge(TbClock);
      end if;
      FT2232H_FSDO <= '0';
      --запись 8 значащих бит
      write8bit : for i in 0 to 7 loop
        wait until rising_edge(TbClock);
        --FT2232H_FSDO <= FullHeader(i + k*8);
        FT2232H_FSDO <= FullHeader(47 - (k * 8 + i));--записываемый бит
      end loop write8bit;
      -- запись Source bit
      wait until rising_edge(TbClock);
      FT2232H_FSDO <= '1';
    end loop full_write;

  end procedure ReadCommand;

begin
  TbClock <= not TbClock after TbPeriod/2 when TbSimEnded /= '1' else '0';
  tester_clk <= TbClock;
  
  
  --установка FT2232H_FSCTS по запросу FT2232H_FSDI на 10 тактов
  set_FT2232H_FSCTS : process(TbClock)
  begin
    if(rising_edge(TbClock)) then
	   if (CTS_open_r = '0' and FT2232H_FSDI = '0') then
		      FSDI_count <= "0000";
	         CTS_open_r <= '1';
				FT2232H_FSCTS <= '0';
		else
				FSDI_count <= std_logic_vector(to_unsigned(to_integer(unsigned(FSDI_count)) + 1, 4));
	   end if;
	 
	   if (CTS_open_r = '1' and FSDI_count = "1000") then 
	       FT2232H_FSCTS <= '1';
	  	    CTS_open_r <= '0';
	   end if;
	 end if;
  end process;

  
  stimuli : process
  begin
    tester_reset <= '0';
    wait for TbPeriod;
    tester_reset <= '1';
    wait for TbPeriod;
	--0000
  --   test_FullHeader <= Test_Concatination("0000000001", '0', "010", TID_count, "0000000100000000");
     WriteCommand("0000000010", '1', "010", TID_count, "0000000000000000", "0100000011111111", FT2232H_FSDO);
	  TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 
	 
	 --read
	--  test_FullHeader <= Test_Concatination("0000000001", '1', "001", TID_count, "0000000100000001");
     ReadCommand("0000000010", '1', "001", TID_count, "0000000000000000", FT2232H_FSDO);
     TID_count <= RecalculationTID(TID_count);
	 
     wait for TbPeriod;
    --0004
	--   test_FullHeader <= Test_Concatination("0000000001", '0', "010", TID_count, "0000000100000000");
     WriteCommand("0000000100", '1', "110", TID_count, "0000001000000100", "00000010001111110000000011111111", FT2232H_FSDO);
	  TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 
	 
	 --101
	--  test_FullHeader <= Test_Concatination("0000000001", '1', "001", TID_count, "0000000100000001");
     ReadCommand("0000000100", '1', "101", TID_count, "0000001000000100", FT2232H_FSDO);
     TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	--0008
	--   test_FullHeader <= Test_Concatination("0000000001", '0', "010", TID_count, "0000000100000000");
     WriteCommand("0000000100", '1', "110", TID_count, "0000001000001000", "00000001000000100000100100100100", FT2232H_FSDO);
	  TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 
	 
	 --101
	--  test_FullHeader <= Test_Concatination("0000000001", '1', "001", TID_count, "0000000100000001");
     ReadCommand("0000000100", '1', "101", TID_count, "0000001000001000", FT2232H_FSDO);
     TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 --000C
	 --   test_FullHeader <= Test_Concatination("0000000001", '0', "010", TID_count, "0000000100000000");
     WriteCommand("0000000010", '1', "110", TID_count, "0000001000001100", "0000000100111110", FT2232H_FSDO);
	  TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 
	 
	 --101
	--  test_FullHeader <= Test_Concatination("0000000001", '1', "001", TID_count, "0000000100000001");
     ReadCommand("0000000010", '1', "101", TID_count, "0000001000001100", FT2232H_FSDO);
     TID_count <= RecalculationTID(TID_count);
     wait for TbPeriod;
	 
	 --CTI
	counter: for k in 0 to 8 loop
		WriteCommand("0011110010", '1', "100", TID_count, "0000001000001100", "000001101001010001010100011000110101111001111000101110111010111000100001000101111011111001010001010100010111101101010111111100110101011110001001001011010001101010000100101011100101001011001101111001100010101000110111110010010001100101101100100001111110001110110111001101011101011011111001101001001100110101011001100110100111110100100101010101010001001100001011000000100010111011000101000000110001010101101010110110100100111111111110111010001000011110001101010011000110011010101011101010010110001101110100011100101001010111010110100111001011101010111111010010111110101100010010111011101001101110100000100001100001101011011000001001100001100000100001000111110101101101101001110000100100001111101101000010111010100000101010010000111000010000000001101111110111110101110011101010000101110111011101111011010011100000011011111100111100001110011110000101100110111000010001100100111001000010110001011111010111100110011110101001000011001000101000011001000110110101000001100111110100000011101010001100110011010000111000101000011100000110110101100111001011000100100010000011110110000000100010010010011111110110011101000110011100000011011010110000110101110101100011000001111001100111011110010101111001011110111111101000111011100011101001111110001000111100000101101101001000110100100111001000100011100110100111000111010010010100011100101100100001111011010110111111010111001011101001111101111110011000000100100000011111100000110000101100001010110110101111110100111110001110101110000001100011011010100101100110001010000111011100011110100001000110111010011110010001111011111101001101011100001110110011011100011001000000010100111111111111100110000111110000100001000011010010100101000111001110010101000100001001000001010101110100011101000011101001110010110101010011011111000010011011100101000011111010100001010111110111000001100101000001010001100110100000010111001011011101100001101100010001101010101011010011010101100101101000011011111010111110011000010010010011111001010001001011110110000001001000010110000110100010101111100001110110001110111010000000000110010111111011110011101011110101100111011001000010100001001011101110010100010100000101011100011111011101101000010000101010010001101011111101111000111000110101110111100000110100000111101011010011001101101001000001001001010110100001001001000100001010101111011101010001001110010001101100100110001100110111011011010001001000110101100101010101111101111010101010010100010110100111100111110101001010101110111010010001011010011000110111101001110000000001001111100111010111100110010001111101101111010100001000011010000001011111011110101111011001101110101010101111010011101111111111101011010010000000101111000011101110011101110010000000101010010001000100001101010100010011001110100110001111000010101000011101101010101000110101000001111000110100111001010101010010100000011111001011011100101000110110101010100010010011010010000111101000011111101000010001111011101011101100010010010000100100111110110101011001111101110100110100011101101110110000001100001101000101001100101000010111100000010000011110110011010000111011000111100000111001111011001011010010101110101001111111100001011101001111000111011111001000011111110000110010001100110100101010110011000111011011010110100001001000011001010000100110010001011101100111111001101100001000010111101000000110011010100101110101101001110101101001100100011111010100001010011001000100000111100110111010110100000010100110100111011011110100010110111101011011001100001001111011101100011011110110010000000110111000101101011000010001110001000000011011011111101001111011011101010011101100101000101010111110011001010011111010111100100100100010110001010101110000100010101000110110111011101100110010000100000101101110110100001111110000010100010111001101110110100011111110001001000111011010101000010001000010111000100101010010101010100001110000010000100111001000100101000000100100110110010101111110100010011111010011000111011100100111000001111001110110111011001010000101110011101001010101001111010110000000011001101110001010100001100110100010010001100001010110011011000001010000100010011100010010001110111101000011111111100111101010010101111110010010000000101000001101100101000001010011001001001000111000011111000010011101101000011010001010011011001101011101100100010011100000001101001101100000000110101011001100011100101001011011000101000100001100010110100000000000110010001111001110001001011111101110001001110000110110001101100010111100110111011110001101101101110110010011111101001101010001010001101111001111001100110101101001101001010011000111100000101110010000111100001010100011101110100000101011110100001101101101101100010000110010101111011011011011111001100010011101110010001110101000111000101111001110110010000101010010110011100101011000010000000001011100001010000100011100100101010100110001100101110101110001011110111101000011111111001010111111001001111000010110110110001010110011010000000000010001110001011011111000111101011100100100001111101101110100001000010011010110000110010011100010001001000001011100111111001000111001110001100110101010110010101101111110101011111001110101101000001110101001110111101101110100110110100100111100000000001100100000100100100011101000101111000001000100011101110010101111010010010011010011101110100111111110001111111100100001111000110111100111100010100110101100100110010111001101110001000111010110001001001001000111000010011000010000111000001011000101100001111011000101011110110101011001000011010000101111101100110001110000100101110000110010010000101011101001011111100010100100000101011110110001000111111100011011000010101110011110100110010100100011110111001110111000110100000101011000110110011101000000101100011101010000111011000101011101001111100100010111010111101001001011011111001000100001110010010100000110101110010100001111110110100010110010011000111010100010011000001101111101101001110010001001001110011000111111000011001000001010001100001010101110000101100111001100001110000100000001000100010010011000100111111001001000011001001100000100011001100011001011111100100010111110010111110100110110110110111011110111000011110001101010000100110101011001011110010101101100100000001111111011011010011000010110000011010101101010110001100110111001101000010111101101101110110100001111001110100101000000000110000010111100000010011011001100110011111001100100011111111011011111101000111100010110111000100111001011011000100110011001001100101111001100010001110001000110010100100011110010111110000000000110011011111101011101111000101000010111010010110000101001111101000111110101000101011100010111101010100100100100100010111110100100000001110100101110100111001001101111011001000011100101110010100100001111101100000011110010000010011001001010011010100100001010111101101001101011110100000100000001001110000100110101101111000000111000000000000111010001110011111011000100101010101110110100011100001011100001101101101010101010111010000111101011010100101001010100010000001100100111011000001100001110000111011010110010000010110100100101101101000110001001010001100110111100100110111011000111110010011101000011000000010100111011001001101100100111011010110001010000000101011011100000111100111001100100110011000001100000010011011111000011001000011111111000111000111110010111000001010010001010011111111001011111010010011111010010010110011000000111011010010010000101010011010110100101100000101010011111000010000010010011110110100011101110100110100000010000001010111001100111110100110011001011101100001010110110100010011101100101001100001110100010010010011111000110101101111010101111001111110101001000101100111101110101110010010100111010101001001101011111101011001110111111000101100001111110011001001100111100011010110111001101111101011110000011000100101000000011111001001100100101101000101010011010000100011010111000001011000000101010010001110101011111101011001100001000100010010010111011010100100010000101011101001000111111100111011000101000011101010011010110011100001100110100111010111100001101010111011011111111011100001110001100110111001001101011100001011011010000000010000000111111101001000101000111110011010011111101011101010000011011000001100101001000110001100000001010110111100001110001011111011101000101011111010001001010110100100010011110001100001011100010000111000010100110010010011010110101000010110100000001101001010001010100011000110101111001111000101110111010111000100001000101111011111001010001010100010111101101010111111100110101011110001001001011010001101010000100101011100101001011001101111001100010101000110111110010010001100101101100100001111110001110110111001101011101011011111001101001001100110101011001100110100111110100100101010101010001001100001011000000100010111011000101000000110001010101101010110110100100111111111110111010001000011110001101010011000110011010101011101010010110001101110100011100101001010111010110100111001011101010111111010010111110101100010010111011101001101110100000100001100001101011011000001001100001100000100001000111110101101101101001110000100100001111101101000010111010100000101010010000111000010000000001101111110111110101110011101010000101110111011101111011010011100000011011111100111100001110011110000101100110111000010001100100111001000010110001011111010111100110011110101001000011001000101000011001000110110101000001100111110100000011101010001100110011010000111000101000011100000110110101100111001011000100100010000011110110000000100010010010011111110110011101000110011100000011011010110000110101110101100011000001111001100111011110010101111001011110111111101000111011100011101001111110001000111100000101101101001000110100100111001000100011100110100111000111010010010100011100101100100001111011010110111111010111001011101001111101111110011000000100100000011111100000110000101100001010110110101111110100111110001110101110000001100011011010100101100110001010000111011100011110100001000110111010011110010001111011111101001101011100001110110011011100011001000000010100111111111111100110000111110000100001000011010010100101000111001110010101000100001001000001010101110100011101000011101001110010110101010011011111000010011011100101000011111010100001010111110111000001100101000001010001100110100000010111001011011101100001101100010001101010101011010011010101100101101000011011111010111110011000010010010011111001010001001011110110000001001000010110000110100010101111100001110110001110111010000000000110010111111011110011101011110101100111011001000010100001001011101110010100010100000101011100011111011101101000010000101010010001101011111101111000111000110101110111100000110100000111101011010011001101101001000001001001010110100001001001000100001010101111011101010001001110010001101100100110001100110111011011010001001000110101100101010101111101111010101010010100010110100111100111110101001010101110111010010001011010011000110111101001110000000001001111100111010111100110010001111101101111010100001000011010000001011111011110101111011001101110101010101111010011101111111111101011010010000000101111000011101110011101110010000000101010010001000100001101010100010011001110100110001111000010101000011101101010101000110101000001111000110100111001010101010010100000011111001011011100101000110110101010100010010011010010000111101000011111101000010001111011101011101100010010010000100100111110110101011001111101110100110100011101101110110000001100001101000101001100101000010111100000010000011110110011010000111011000111100000111001111011001011010010101110101001111111100001011101001111000111011111001000011111110000110010001100110100101010110011000111011011010110100001001000011001010000100110010001011101100111111001101100001000010111101000000110011010100101110101101001110101101001100100011111010100001010011001000100000111100110111010110100000010100110100111011011110100010110111101011011001100001001111011101100011011110110010000000110111000101101011000010001110001000000011011011111101001111011011101010011101100101000101010111110011001010011111010111100100100100010110001010101110000100010101000110110111011101100110010000100000101101110110100001111110000010100010111001101110110100011111110001001000111011010101000010001000010111000100101010010101010100001110000010000100111001000100101000000100100110110010101111110100010011111010011000111011100100111000001111001110110111011001010000101110011101001010101001111010110000000011001101110001010100001100110100010010001100001010110011011000001010000100010011100010010001110111101000011111111100111101010010101111110010010000000101000001101100101000001010011001001001000111000011111000010011101101000011010001010011011001101011101100100010011100000001101001101100000000110101011001100011100101001011011000101000100001100010110100000000000110010001111001110001001011111101110001001110000110110001101100010111100110111011110001101101101110110010011111101001101010001010001101111001111001100110101101001101001010011000111100000101110010000111100001010100011101110100000101011110100001101101101101100010000110010101111011011011011111001100010011101110010001110101000111000101111001110110010000101010010110011100101011000010000000001011100001010000100011100100101010100110001100101110101110001011110111101000011111111001010111111001001111000010110110110001010110011010000000000010001110001011011111000111101011100100100001111101101110100001000010011010110000110010011100010001001000001011100111111001000111001110001100110101010110010101101111110101011111001110101101000001110101001110111101101110100110110100100111100000000001100100000100100100011101000101111000001000100011101110010101111010010010011010011101110100111111110001111111100100001111000110111100111100010100110101100100110010111001101110001000111010110001001001001000111000010011000010000111000001011000101100001111011000101011110110101011001000011010000101111101100110001110000100101110000110010010000101011101001011111100010100100000101011110110001000111111100011011000010101110011110100110010100100011110111001110111000110100000101011000110110011101000000101100011101010000111011000101011101001111100100010111010111101001001011011111001000100001110010010100000110101110010100001111110110100010110010011000111010100010011000001101111101101001110010001001001110011000111111000011001000001010001100001010101110000101100111001100001110000100000001000100010010011000100111111001001000011001001100000100011001100011001011111100100010111110010111110100110110110110111011110111000011110001101010000100110101011001011110010101101100100000001111111011011010011000010110000011010101101010110001100110111001101000010111101101101110110100001111001110100101000000000110000010111100000010011011001100110011111001100100011111111011011111101000111100010110111000100111001011011000100110011001001100101111001100010001110001000110010100100011110010111110000000000110011011111101011101111000101000010111010010110000101001111101000111110101000101011100010111101010100100100100100010111110100100000001110100101110100111001001101111011001000011100101110010100100001111101100000011110010000010011001001010011010100100001010111101101001101011110100000100000001001110000100110101101111000000111000000000000111010001110011111011000100101010101110110100011100001011100001101101101010101010111010000111101011010100101001010100010000001100100111011000001100001110000111011010110010000010110100100101101101000110001001010001100110111100100110111011000111110010011101000011000000010100111011001001101100100111011010110001010000000101011011100000111100111001100100110011000001100000010011011111000011001000011111111000111000111110010111000001010010001010011111111001011111010010011111010010010110011000000111011010010010000101010011010110100101100000101010011111000010000010010011110110100011101110100110100000010000001010111001100111110100110011001011101100001010110110100010011101100101001100001110100010010010011111000110101101111010101111001111110101001000101100111101110101110010010100111010101001001101011111101011001110111111000101100001111110011001001100111100011010110111001101111101011110000011000100101000000011111001001100100101101000101010011010000100011010111000001011000000101010010001110101011111101011001100001000100010010010111011010100100010000101011101001000111111100111011000101000011101010011010110011100001100110100111010111100001101010111011011111111011100001110001100110111001001101011100001011011010000000010000000111111101001000101000111110011010011111101011101010000011011000001100101001000110001100000001010110111100001110001011111011101000101011111010001001010110100100010011110001100001011100010000111000010100110010010011010110101000010110100000001101001010001010100011000110101111001111000101110111010111000100001000101111011111001010001010100010111101101010111111100110101011110001001001011010001101010000100101011100101001011001101111001100010101000110111110010010001100101101100100001111110001110110111001101011101011011111001101001001100110101011001100110100111110100100101010101010001001100001011000000100010111011000101000000110001010101101010110110100100111111111110111010001000011110001101010011000110011010101011101010010110001101110100011100101001010111010110100111001011101010111111010010111110101100010010111011101001101110100000100001100001101011011000001001100001100000100001000111110101101101101001110000100100001111101101000010111010100000101010010000111000010000000001101111110111110101110011101010000101110111011101111011010011100000011011111100111100001110011110000101100110111000010001100100111001000010110001011111010111100110011110101001000011001000101000011001000110110101000001100111110100000011101010001100110011010000111000101000011100000110110101100111001011000100100010000011110110000000100010010010011111110110011101000110011100000011011010110000110101110101100011000001111001100111011110010101111001011110111111101000111011100011101001111110001000111100000101101101001000110100100111001000100011100110100111000111010010010100011100101100100001111011010110111111010111001011101001111101111110011000000100100000011111100000110000101100001010110110101111110100111110001110101110000001100011011010100101100110001010000111011100011110100001000110111010011110010001111011111101001101011100001110110011011100011001000000010100111111111111100110000111110000100001000011010010100101000111001110010101000100001001000001010101110100011101000011101001110010110101010011011111000010011011100101000011111010100001010111110111000001100101000001010001100110100000010111001011011101100001101100010001101010101011010011010101100101101000011011111010111110011000010010010011111001010001001011110110000001001000010110000110100010101111100001110110001110111010000000000110010111111011110011101011110101100111011001000010100001001011101110010100010100000101011100011111011101101000010000101010010001101011111101111000111000110101110111100000110100000111101011010011001101101001000001001001010110100001001001000100001010101111011101010001001110010001101100100110001100110111011011010001001000110101100101010101111101111010101010010100010110100111100111110101001010101110111010010001011010011000110111101001110000000001001111100111010111100110010001111101101111010100001000011010000001011111011110101111011001101110101010101111010011101111111111101011010010000000101111000011101110011101110010000000101010010001000100001101010100010011001110100110001111000010101000011101101010101000110101000001111000110100111001010101010010100000011111001011011100101000110110101010100010010011010010000111101000011111101000010001111011101011101100010010010000100100111110110101011001111101110100110100011101101110110000001100001101000101001100101000010111100000010000011110110011010000111011000111100000111001111011001011010010101110101001111111100001011101001111000111011111001000011111110000110010001100110100101010110011000111011011010110100001001000011001010000100110010001011101100111111001101100001000010111101000000110011010100101110101101001110101101001100100011111010100001010011001000100000111100110111010110100000010100110100111011011110100010110111101011011001100001001111011101100011011110110010000000110111000101101011000010001110001000000011011011111101001111011011101010011101100101000101010111110011001010011111010111100100100100010110001010101110000100010101000110110111011101100110010000100000101101110110100001111110000010100010111001101110110100011111110001001000111011010101000010001000010111000100101010010101010100001110000010000100111001000100101000000100100110110010101111110100010011111010011000111011100100111000001111001110110111011001010000101110011101001010101001111010110000000011001101110001010100001100110100010010001100001010110011011000001010000100010011100010010001110111101000011111111100111101010010101111110010010000000101000001101100101000001010011001001001000111000011111000010011101101000011010001010011011001101011101100100010011100000001101001101100000000110101011001100011100101001011011000101000100001100010110100000000000110010001111001110001001011111101110001001110000110110001101100010111100110111011110001101101101110110010011111101001101010001010001101111001111001100110101101001101001010011000111100000101110010000111100001010100011101110100000101011110100001101101101101100010000110010101111011011011011111001100010011101110010001110101000111000101111001110110010000101010010110011100101011000010000000001011100001010000100011100100101010100110001100101110101110001011110111101000011111111001010111111001001111000010110110110001010110011010000000000010001110001011011111000111101011100100100001111101101110100001000010011010110000110010011100010001001000001011100111111001000111001110001100110101010110010101101111110101011111001110101101000001110101001110111101101110100110110100100111100000000001100100000100100100011101000101111000001000100011101110010101111010010010011010011101110100111111110001111111100100001111000110111100111100010100110101100100110010111001101110001000111010110001001001001000111000010011000010000111000001011000101100001111011000101011110110101011001000011010000101111101100110001110000100101110000110010010000101011101001011111100010100100000101011110110001000111111100011011000010101110011110100110010100100011110111001110111000110100000101011000110110011101000000101100011101010000111011000101011101001111100100010111010111101001001011011111001000100001110010010100000110101110010100001111110110100010110010011000111010100010011000001101111101101001110010001001001110011000111111000011001000001010001100001010101110000101100111001100001110000100000001000100010010011000100111111001001000011001001100000100011001100011001011111100100010111110010111110100110110110110111011110111000011110001101010000100110101011001011110010101101100100000001111111011011010011000010110000011010101101010110001100110111001101000010111101101101110110100001111001110100101000000000110000010111100000010011011001100110011111001100100011111111011011111101000111100010110111000100111001011011000100110011001001100101111001100010001110001000110010100100011110010111110000000000110011011111101011101111000101000010111010010110000101001111101000111110101000101011100010111101010100100100100100010111110100100000001110100101110100111001001101111011001000011100101110010100100001111101100000011110010000010011001001010011010100100001010111101101001101011110100000100000001001110000100110101101111000000111000000000000111010001110011111011000100101010101110110100011100001011100001101101101010101010111010000111101011010100101001010100010000001100100111011000001100001110000111011010110010000010110100100101101101000110001001010001100110111100100110111011000111110010011101000011000000010100111011001001101100100111011010110001010000000101011011100000111100111001100100110011000001100000010011011111000011001000011111111000111000111110010111000001010010001010011111111001011111010010011111010010010110011000000111011010010010000101010011010110100101100000101010011111000010000010010011110110100011101110100110100000010000001010111001100111110100110011001011101100001010110110100010011101100101001100001110100010010010011111000110101101111010101111001111110101001000101100111101110101110010010100111010101001001101011111101011001110111111000101100001111110011001001100111100011010110111001101111101011110000011000100101000000011111001001100100101101000101010011010000100011010111000001011000000101010010001110101011111101011001100001000100010010010111011010100100010000101011101001000111111100111011000101000011101010011010110011100001100110100111010111100001101010111011011111111011100001110001100110111001001101011100001011011010000000010000000111111101001000101000111110011010011111101011101010000011011000001100101001000110001100000001010110111100001110001011111011101000101011111010001001010110100100010011110001100001011100010000111000010100110010010011010110101000010110100000001101001010001010100011000110101111001111000101110111010111000100001000101111011111001010001010100010111101101010111111100110101011110001001001011010001101010000100101011100101001011001101111001100010101000110111110010010001100101101100100001111110001110110111001101011101011011111001101001001100110101011001100110100111110100100101010101010001001100001011000000100010111011000101000000110001010101101010110110100100111111111110111010001000011110001101010011000110011010101011101010010110001101110100011100101001010111010110100111001011101010111111010010111110101100010010111011101001101110100000100001100001101011011000001001100001100000100001000111110101101101101001110000100100001111101101000010111010100000101010010000111000010000000001101111110111110101110011101010000101110111011101111011010011100000011011111100111100001110011110000101100110111000010001100100111001000010110001011111010111100110011110101001000011001000101000011001000110110101000001100111110100000011101010001100110011010000111000101000011100000110110101100111001011000100100010000011110110000000100010010010011111110110011101000110011100000011011010110000110101110101100011000001111001100111011110010101111001011110111111101000111011100011101001111110001000111100000101101101001000110100100111001000100011100110100111000111010010010100011100101100100001111011010110111111010111001011101001111101111110011000000100100000011111100000110000101100001010110110101111110100111110001110101110000001100011011010100101100110001010000111011100011110100001000110111010011110010001111011111101001101011100001110110011011100011001000000010100111111111111100110000111110000100001000011010010100101000111001110010101000100001001000001010101110100011101000011101001110010110101010011011111000010011011100101000011111010100001010111110111000001100101000001010001100110100000010111001011011101100001101100010001101010101011010011010101100101101000011011111010111110011000010010010011111001010001001011110110000001001000010110000110100010101111100001110110001110111010000000000110010111111011110011101011110101100111011001000010100001001011101110010100010100000101011100011111011101101000010000101010010001101011111101111000111000110101110111100000110100000111101011010011001101101001000001001001010110100001001001000100001010101111011101010001001110010001101100100110001100110111011011010001001000110101100101010101111101111010101010010100010110100111100111110101001010101110111010010001011010011000110111101001110000000001001111100111010111100110010001111101101111010100001000011010000001011111011110101111011001101110101010101111010011101111111111101011010010000000101111000011101110011101110010000000101010010001000100001101010100010011001110100110001111000010101000011101101010101000110101000001111000110100111001010101010010100000011111001011011100101000110110101010100010010011010010000111101000011111101000010001111011101011101100010010010000100100111110110101011001111101110100110100011101101110110000001100001101000101001100101000010111100000010000011110110011010000111011000111100000111001111011001011010010101110101001111111100001011101001111000111011111001000011111110000110010001100110100101010110011000111011011010110100001001000011001010000100110010001011101100111111001101100001000010111101000000110011010100101110101101001110101101001100100011111010100001010011001000100000111100110111010110100000010100110100111011011110100010110111101011011001100001001111011101100011011110110010000000110111000101101011000010001110001000000011011011111101001111011011101010011101100101000101010111110011001010011111010111100100100100010110001010101110000100010101000110110111011101100110010000100000101101110110100001111110000010100010111001101110110100011111110001001000111011010101000010001000010111000100101010010101010100001110000010000100111001000100101000000100100110110010101111110100010011111010011000111011100100111000001111001110110111011001010000101110011101001010101001111010110000000011001101110001010100001100110100010010001100001010110011011000001010000100010011100010010001110111101000011111111100111101010010101111110010010000000101000001101100101000001010011001001001000111000011111000010011101101000011010001010011011001101011101100100010011100000001101001101100000000110101011001100011100101001011011000101000100001100010110100000000000110010001111001110001001011111101110001001110000110110001101100010111100110111011110001101101101110110010011111101001101010001010001101111001111001100110101101001101001010011000111100000101110010000111100001010100011101110100000101011110100001101101101101100010000110010101111011011011011111001100010011101110010001110101000111000101111001110110010000101010010110011100101011000010000000001011100001010000100011100100101010100110001100101110101110001011110111101000011111111001010111111001001111000010110110110001010110011010000000000010001110001011011111000111101011100100100001111101101110100001000010011010110000110010011100010001001000001011100111111001000111001110001100110101010110010101101111110101011111001110101101000001110101001110111101101110100110110100100111100000000001100100000100100100011101000101111000001000100011101110010101111010010010011010011101110100111111110001111111100100001111000110111100111100010100110101100100110010111001101110001000111010110001001001001000111000010011000010000111000001011000101100001111011000101011110110101011001000011010000101111101100110001110000100101110000110010010000101011101001011111100010100100000101011110110001000111111100011011000010101110011110100110010100100011110111001110111000110100000101011000110110011101000000101100011101010000111011000101011101001111100100010111010111101001001011011111001000100001110010010100000110101110010100001111110110100010110010011000111010100010011000001101111101101001110010001001001110011000111111000011001000001010001100001010101110000101100111001100001110000100000001000100010010011000100111111001001000011001001100000100011001100011001011111100100010111110010111110100110110110110111011110111000011110001101010000100110101011001011110010101101100100000001111111011011010011000010110000011010101101010110001100110111001101000010111101101101110110100001111001110100101000000000110000010111100000010011011001100110011111001100100011111111011011111101000111100010110111000100111001011011000100110011001001100101111001100010001110001000110010100100011110010111110000000000110011011111101011101111000101000010111010010110000101001111101000111110101000101011100010111101010100100100100100010111110100100000001110100101110100111001001101111011001000011100101110010100100001111101100000011110010000010011001001010011010100100001010111101101001101011110100000100000001001110000100110101101111000000111000000000000111010001110011111011000100101010101110110100011100001011100001101101101010101010111010000111101011010100101001010100010000001100100111011000001100001110000111011010110010000010110100100101101101000110001001010001100110111100100110111011000111110010011101000011000000010100111011001001101100100111011010110001010000000101011011100000111100111001100100110011000001100000010011011111000011001000011111111000111000111110010111000001010010001010011111111001011111010010011111010010010110011000000111011010010010000101010011010110100101100000101010011111000010000010010011110110100011101110100110100000010000001010111001100111110100110011001011101100001010110110100010011101100101001100001110100010010010011111000110101101111010101111001111110101001000101100111101110101110010010100111010101001001101011111101011001110111111000101100001111110011001001100111100011010110111001101111101011110000011000100101000000011111001001100100101101000101010011010000100011010111000001011000000101010010001110101011111101011001100001000100010010010111011010100100010000101011101001000111111100111011000101000011101010011010110011100001100110100111010111100001101010111011011111111011100001110001100110111001001101011100001011011010000000010000000111111101001000101000111110011010011111101011101010000011011000001100101001000110001100000001010110111100001110001011111011101000101011111010001001010110100100010011110001100001011100010000111000010100110010010011010110101000010110100", FT2232H_FSDO);
		TID_count <= RecalculationTID(TID_count);
		wait for TbPeriod;
	end loop counter ;
	skiptime(10);
	wait for TbPeriod;
	read_counter: for k in 0 to 10 loop
		 ReadCommand("0011110010", '1', "011", TID_count, "0000001000001100", FT2232H_FSDO);
		 TID_count <= RecalculationTID(TID_count);
		 wait for TbPeriod;
	end loop read_counter ;
    skiptime(3000);
    TbSimEnded <= '1';
  end process;
  

end tester_top;
configuration ts_top of Tester is
  for tester_top
  end for;
end ts_top;